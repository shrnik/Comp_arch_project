`timescale 1ns/10ps
module mux_16x1(y,a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,s);
input [n-1:0]a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15;
input [3:0]s;
output reg [n-1:0]y;
parameter n = 16;

always @(*)
begin
case (s)
4'b0000: y=a0;
4'b0001: y=a1;
4'b0010: y=a2;
4'b0011: y=a3;
4'b0100: y=a4;
4'b0101: y=a5;
4'b0110: y=a6;
4'b0111: y=a7;
4'b1000: y=a8;
4'b1001: y=a9;
4'b1010: y=a10;
4'b1011: y=a11;
4'b1100: y=a12;
4'b1101: y=a13;
4'b1110: y=a14;
4'b1111: y=a15;
endcase
end
endmodule
module tb_mux_16x1();
wire [n-1:0]y;
reg [n-1:0]a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15;
reg [3:0]s;
parameter n=16;

mux_16x1 uut(y,a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,s);
initial $monitor("t=%3d, y=%16b, a0=%16b, a1=%16b, a2=%16b, a3=%16b, a4=%16b, a5=%16b, a6=%16b, a7=%16b, a8=%16b, a9=%16b, a10=%16b, a11=%16b, a12=%16b, a13=%16b, a14=%16b, a15=%16b,  s=%4b",$time,y,a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,s);
initial     
	begin      
$dumpfile("mux_16x1.vcd");    
$dumpvars;     
end 

initial
	begin 
		#010 a0  = 16'b1111111111111110 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#010 s = 4'b0000;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111101 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b0001;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111011 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b0010;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111110111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b0011;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b0100;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b0101;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b0110;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b0111;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1000;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1001;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1010;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1011;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1100;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1101;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1110;
		#010 a0  = 16'b1111111111111111 ; a1  = 16'b1111111111111111 ; a2  = 16'b1111111111111111 ; a3  = 16'b1111111111111111 ; a4  = 16'b1111111111111111 ; a5  = 16'b1111111111111111 ; a6  = 16'b1111111111111111 ; a7  = 16'b1111111111111111 ; a8  = 16'b1111111111111111 ; a9  = 16'b1111111111111111 ; a10  = 16'b1111111111111111 ; a11  = 16'b1111111111111111 ; a12  = 16'b1111111111111111 ; a13  = 16'b1111111111111111 ; a14  = 16'b1111111111111111 ; a15  = 16'b1111111111111111 ; 
		#020 s = 4'b1111;
		end
initial 
#1000 $stop;
endmodule
		