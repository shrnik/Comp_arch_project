`timescale 1ns/10ps
module dec_4x16(a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,s);
output reg a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15;
input [3:0]s;

always @ (s)
begin
a0=1'b0;  a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0;

	case(s)
	4'b0000: a0=1'b1;/*   a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b0001: a1=1'b1;  /* a1=1'b1; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b0010: a2=1'b1;  /* a1=1'b0; a2=1'b1; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b0011: a3=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b1; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b0100: a4=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b1; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b0101: a5=1'b1; /*  a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b1; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b0110: a6=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b1; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b0111: a7=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b1; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b1000: a8=1'b1; /*  a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b1; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b1001: a9=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b1; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b1010: a10=1'b1; /*  a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b1; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b1011: a11=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b1; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b1100: a12=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b1; a13=1'b0; a14=1'b0;  a15=1'b0; */
	4'b1101: a13=1'b1;  /* a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b1; a14=1'b0;  a15=1'b0; */
	4'b1110: a14=1'b1; /*  a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b1;  a15=1'b0; */
	4'b1111: a15=1'b1; /*  a1=1'b0; a2=1'b0; a3=1'b0; a4=1'b0; a5=1'b0; a6=1'b0; a7=1'b0; a8=1'b0; a9=1'b0; a10=1'b0; a11=1'b0; a12=1'b0; a13=1'b0; a14=1'b0;  a15=1'b1; */
	endcase
	end
endmodule	

module tb_dec_4x16();
wire a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15;
reg [3:0]s;

dec_4x16 uut(a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,s);
initial $monitor("t=%3d, a0=%1b, a1=%1b, a2=%1b, a3=%1b, a4=%1b, a5=%1b, a6=%1b, a7=%1b, a8=%1b, a9=%1b, a10=%1b, a11=%1b, a12=%1b, a13=%1b, a14=%1b, a15=%1b,  s=%4b",$time,a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,s);
initial     
	begin      
$dumpfile("dec_4x16.vcd");    
$dumpvars;     
end 

initial
	begin 
		#010 s = 4'b0000;
		#020 s = 4'b0001;
		#020 s = 4'b0010;
		#020 s = 4'b0011;
		#020 s = 4'b0100;
		#020 s = 4'b0101;
		#020 s = 4'b0110;
		#020 s = 4'b0111;
		#020 s = 4'b1000;
		#020 s = 4'b1001;
		#020 s = 4'b1010;
		#020 s = 4'b1011;
		#020 s = 4'b1100;
		#020 s = 4'b1101;
		#020 s = 4'b1110;
		#020 s = 4'b1111;
		end
initial 
#1000 $stop;
endmodule